// I worked on building a circuit to process scancodes from a PS/2 keyboard for a game. The challenge involved recognizing specific scancodes for arrow keys and asserting the correct output using a case statement.


module top_module (
    input [15:0] scancode,
    output reg left,
    output reg down,
    output reg right,
    output reg up
);

always @(*) begin
    {up, down, left, right} = 4'b0;
    case (scancode)
        16'he06b: left = 1;
        16'he072: down = 1;
        16'he074: right = 1;
        16'he075: up = 1;
    endcase
end

endmodule
